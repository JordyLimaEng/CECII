module decoder(input logic [4:0] a,
 output logic [31:0] y);
 
 always_comb
 case(a)
 5'd00: y = 32'b00000000000000000000000000000000;
 5'd01: y = 32'b00000000000000000000000000000001;
 5'd02: y = 32'b00000000000000000000000000000010;
 5'd03: y = 32'b00000000000000000000000000000100;
 5'd04: y = 32'b00000000000000000000000000001000;
 5'd05: y = 32'b00000000000000000000000000010000;
 5'd06: y = 32'b00000000000000000000000000100000;
 5'd07: y = 32'b00000000000000000000000001000000;
 5'd08: y = 32'b00000000000000000000000010000000;
 5'd09: y = 32'b00000000000000000000000100000000;
 5'd10: y = 32'b00000000000000000000001000000000;
 5'd11: y = 32'b00000000000000000000010000000000;
 5'd12: y = 32'b00000000000000000000100000000000;
 5'd13: y = 32'b00000000000000000001000000000000;
 5'd14: y = 32'b00000000000000000010000000000000;
 5'd15: y = 32'b00000000000000001000000000000000;
 5'd16: y = 32'b00000000000000010000000000000000;
 5'd17: y = 32'b00000000000000100000000000000000;
 5'd18: y = 32'b00000000000001000000000000000000;
 5'd19: y = 32'b00000000000010000000000000000000;
 5'd20: y = 32'b00000000000100000000000000000000;
 5'd21: y = 32'b00000000001000000000000000000000;
 5'd22: y = 32'b00000000010000000000000000000000;
 5'd23: y = 32'b00000000100000000000000000000000;
 5'd24: y = 32'b00000001000000000000000000000000;
 5'd25: y = 32'b00000010000000000000000000000000;
 5'd26: y = 32'b00000100000000000000000000000000;
 5'd27: y = 32'b00001000000000000000000000000000;
 5'd28: y = 32'b00010000000000000000000000000000;
 5'd29: y = 32'b00100000000000000000000000000000;
 5'd30: y = 32'b01000000000000000000000000000000;
 5'd31: y = 32'b10000000000000000000000000000000;
 default: y=32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
 endcase
 endmodule
 
 