0_0000_Z
0_1111_Z
1_0000_0000
1_1111_1111
