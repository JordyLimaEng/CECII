0_0000_ZZZZ
0_1111_ZZZZ
1_0000_0000
1_1111_1111
